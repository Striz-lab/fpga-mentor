module clk_div(
/*
*   describe ports here
*/
);

/*
*   describe X width register
*/

/*
*   write your clock divider logic here
*/

endmodule

module clk_div_cheats(
/*
*   describe ports here
*/
);

/*
*   paste .veo code here
*/

endmodule