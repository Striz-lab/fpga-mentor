module weird_logic(
/*
*   Problem 1/5:
*   describe ports here
*/
);

/*
*   Problem 1/5:
*   describe your logic here
*/

endmodule