module test(
    input wire in,
    output wire out
);

assign out = in;

endmodule


module invertor(
/*
*   Problem 1/5:
*   describe ports here
*/
);

/*
*   Problem 1/5:
*   write NOT logic here
*/

endmodule